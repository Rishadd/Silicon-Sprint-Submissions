`timescale 1ns / 1ps


module main_decoder();
    // The main decoder interprets the opcode field and produces
    // control signals for the datapath components.    
    
    
endmodule
