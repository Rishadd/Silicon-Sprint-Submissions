`timescale 1ns / 1ps


module single_cycle(clk, rst);

input clk,rst;

    // This is the top-level CPU wrapper - the "brain + body".


    //   Combine all modules built so far into a working single-cycle CPU.
endmodule
