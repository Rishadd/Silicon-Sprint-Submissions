`timescale 1ns / 1ps


module alu_decoder ();
    // The ALU decoder refines control signals. 
    
    // The goal is to produce a 4-bit alu_ctrl that matches the
    // operation encodings used inside your ALU module.
    
    
endmodule
